module IP_tb();

endmodule