
module unsaved (
	clk_clk,
	pio_export,
	reset_reset_n);	

	input		clk_clk;
	inout	[4:0]	pio_export;
	input		reset_reset_n;
endmodule
